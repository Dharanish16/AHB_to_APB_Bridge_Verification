

package test_pkg;

    //import uvm_pkg.sv
	import uvm_pkg::*;

    //include uvm_macros.sv
	`include "uvm_macros.svh"

    `include "ahb_xtn.sv"
    `include "ahb_agt_config.sv"
    `include "apb_agt_config.sv"
    `include "env_config.sv"

    `include "ahb_agt_drv.sv"
    `include "ahb_agt_mon.sv"
    `include "ahb_agt_seqr.sv"
    `include "ahb_agent.sv"
    `include "ahb_agt_top.sv"
    `include "ahb_sequence.sv"

    `include "apb_xtn.sv"
    //`include "normal_seq.sv"
    `include "apb_agt_mon.sv"
    `include "apb_agt_seqr.sv"
    `include "apb_agt_drv.sv"
    `include "apb_agent.sv"
    `include "apb_agt_top.sv"
    

    //`include "virtual_sequencer.sv"
    //`include "virtual_sequence.sv"
    `include "bridge_scoreboard.sv"

    `include "bridge_env.sv"


    `include "ahb2apb_test.sv"

endpackage